
 module mips_16
 endmodule  